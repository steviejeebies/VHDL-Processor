-- Michael Manzke
-- michael.manzke@cs.tcd.ie
-- 25 April 2003

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity control_mem_256x28 is
    Port ( MW : out std_logic;
           MM : out std_logic;
           RW : out std_logic;
           MD : out std_logic;
           FS : out std_logic_vector(4 downto 0);
           MB : out std_logic;
           TB : out std_logic;
           TA : out std_logic;
           TD : out std_logic;
           PL : out std_logic;
           PI : out std_logic;
           IL : out std_logic;
           MC : out std_logic;
           MS : out std_logic_vector(2 downto 0);
           NA : out std_logic_vector(7 downto 0);
           IN_CAR : in std_logic_vector(7 downto 0));
end control_mem_256x28;

architecture behavioural of control_mem_256x28 is
    type mem_array is array (0 to 255) of std_logic_vector(27 downto 0);
    
    begin
        memory_m : process (IN_CAR)
            variable control_mem : mem_array :=(
                                                --0
                                                X"C020224", --0
                                                X"C02000C", --1
                                                X"C020001", --2
                                                X"C020014", --3
                                                X"C0200E4", --4
                                                X"C020024", --5
                                                X"C0E0000", --6     // Branch if Zero Set this instruction checks if the condition NOT Z is true, in which case it continues to C0. Else it increments to the next CAR address
                                                X"C022000", --7     // Branch This instruction has PC load what is in DR and SB, and then also updates CAR to be NA (which points to IF)
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --1
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --2
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --3
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --4
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --5
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --6
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --7
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --8
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --9
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --A
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --B
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --C
                                                X"C10C002", --0
                                                X"0030000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --D
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --E
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"0000000", --6
                                                X"0000000", --7
                                                X"0000000", --8
                                                X"0000000", --9
                                                X"0000000", --A
                                                X"0000000", --B
                                                X"0000000", --C
                                                X"0000000", --D
                                                X"0000000", --E
                                                X"0000000", --F
                                                --F
                                                X"0000000", --0
                                                X"0000000", --1
                                                X"0000000", --2
                                                X"0000000", --3
                                                X"0000000", --4
                                                X"0000000", --5
                                                X"1024000", --6
                                                X"F624000", --7
                                                X"F724000", --8
                                                X"F824000", --9
                                                X"F924000", --A
                                                X"FA20000", --B
                                                X"FB20000", --C
                                                X"FC20000", --D
                                                X"FD20000", --E
                                                X"FE20000"  --F
                                                );

            variable addr : integer;    -- instantiate address to IF for RESET
            variable control_out : std_logic_vector(27 downto 0);
            
            begin
                addr := conv_integer(IN_CAR);
                control_out := control_mem(addr);
                MW <= control_out(0);
                MM <= control_out(1);
                RW <= control_out(2);
                MD <= control_out(3);
                FS <= control_out(8 downto 4);
                MB <= control_out(9);
                TB <= control_out(10);
                TA <= control_out(11);
                TD <= control_out(12);
                PL <= control_out(13);
                PI <= control_out(14);
                IL <= control_out(15);
                MC <= control_out(16);
                MS <= control_out(19 downto 17);
                NA <= control_out(27 downto 20);
            end process;
end behavioural;
                
                                                          
                                                
                                                
           